`define ALU_OP_ADD	8'd0
`define ALU_OP_SLT	8'd1
`define ALU_OP_SLTU	8'd2
`define ALU_OP_AND	8'd3
`define ALU_OP_OR	8'd4
`define ALU_OP_XOR	8'd5
`define ALU_OP_SLL	8'd6
`define ALU_OP_SRL	8'd7
`define ALU_OP_SUB	8'd8
`define ALU_OP_SRA	8'd9
`define ALU_OP_EQ	8'd10
`define ALU_OP_MUL	8'd11
`define ALU_OP_DIV	8'd12
